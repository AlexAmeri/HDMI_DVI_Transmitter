----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/30/2020 10:17:55 PM
-- Design Name: 
-- Module Name: DVI_Transmitter - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity DVI_Transmitter is
      Port (
            --Clocks
            clk : in std_logic;
      
            --VGA inputs
            r_vga, b_vga : in std_logic_vector(4 downto 0);
            g_vga : in std_logic_vector(5 downto 0);
            h_sync, v_sync : in std_logic;
            
            --Control Signals
            vid : in std_logic;
            
            --Outputs
            hdmi_d_p : out std_logic_vector(2 downto 0);
            hdmi_d_n : out std_logic_vector(2 downto 0);
            hdmi_clk_p : out std_logic;
            hdmi_clk_n : out std_logic;
            hdmi_out_en : out std_logic
            
             );
end DVI_Transmitter;

architecture Behavioral of DVI_Transmitter is

    --Components
    --TDMS Encoders
    component tdmi_transmitter is
    Port ( --Control signals shared with VGA logic
           clk, en : in STD_LOGIC;
           
           --HDMI Control signals
           CTL : in std_logic_vector(1 downto 0);
           DE : in std_logic;
           
           --Data input
           dc : in std_logic_vector(7 downto 0);
           
           --Serial Data output
           TDMI_output : out std_logic_vector(9 downto 0)
           );
    end component;    
    
    --Serializer
    component tdms_serializer_combined is
    Port (
        data_red, data_green, data_blue : in std_logic_vector(9 downto 0);
        clk : in std_logic; 
        
        --Blue is 0, Green is 1, Red is 2
        TDMS_out, TDMS_out_not : out std_logic_vector (2 downto 0);
        new_character_clock : out std_logic;
        en : in std_logic
     );
    end component;
  

    --Clock generator
    component DVI_Clock_Generator is
    Port (
        reset : in std_logic;
        base_clk : in std_logic;                --125 MHz base clock
        out_clk_base : out std_logic;           --125 MHz base clock, phase matched to 250 MHz clock
        out_clk_serializer : out std_logic;     --250 MHz serializer clock
        out_clk_en : out std_logic              --25 MHZ clock enable chirp, phase matched to 250 MHz clock
    );
    end component;
    
    --Signals
    --Clocking Signals
    --signal serial_clk : std_logic;
    signal TDMS_character_clock : std_logic;
    signal artificial_base_clk : std_logic;
    signal artificial_clk_en : std_logic;
    signal serializer_bit_clk : std_logic;
    signal r_tdms_bus, g_tdms_bus, b_tdms_bus : std_logic_vector(9 downto 0);
    
    --TDMS Encoder Input Words
    signal r_ctl, g_ctl, b_ctl : std_logic_vector(1 downto 0) := (others => '1');
    
    --TMDS Serializer output data streams
    --Blue is 0, Green is 1, Red is 2
    signal TMDS_stream, TMDS_stream_not : std_logic_vector(2 downto 0);
    
    --FIFO signals
    signal rin, r1, r2, r3, r4 : std_logic_vector(7 downto 0) := (others => '0');
    signal gin, g1, g2, g3, g4 : std_logic_vector(7 downto 0) := (others => '0');
    signal bin, b1, b2, b3, b4 : std_logic_vector(7 downto 0) := (others => '0');
    signal de_in, de1, de2, de3, de4 : std_logic := '0';
    signal hs_in, hs1, hs2, hs3, hs4 : std_logic := '0';
    signal vs_in, vs1, vs2, vs3, vs4 : std_logic := '0';
    
begin

    --Output Buffers, for TMDS
    --Output Differential Signaling Buffers
    OBUFDS_blue  : OBUFDS port map ( O  => hdmi_d_p(0), OB => hdmi_d_n(0), I  => TMDS_stream(0)  );
    OBUFDS_red   : OBUFDS port map ( O  => hdmi_d_p(2), OB => hdmi_d_n(2), I  => TMDS_stream(2) );
    OBUFDS_green : OBUFDS port map ( O  => hdmi_d_p(1), OB => hdmi_d_n(1), I  => TMDS_stream(1)   );
    OBUFDS_clock : OBUFDS port map ( O  => hdmi_clk_p, OB => hdmi_clk_n, I  => TDMS_character_clock );

    --Glue logic
    b_ctl <= vs4 & hs4;
    g_ctl <= "00";
    r_ctl <= "00";
    hdmi_out_en <= '1';
    
    --Make a 5 stage FIFO pipeline for input signals.
    --Since there is a possibility that the DVI clock - generated by an MMCM -
    --is out of phase with the clock used by other user IP, for the sake of robustness
    --a 5 stage FIFO is being used for each input pin.
    rin <= r_vga & "000";
    gin <= g_vga & "00";
    bin <= b_vga & "000";
    de_in <= vid;
    hs_in <= h_sync;
    vs_in <= v_sync;
    
    data_input_pipeline : process(clk)
    begin
        --Advance the FIFO pipeline to prevent clock domain crossing problems
        if(rising_edge(artificial_base_clk)) then
            --Color Signals
            r1 <= rin;
            r2 <= r1;
            r3 <= r2;
            r4 <= r3;
            
            g1 <= gin;
            g2 <= g1;
            g3 <= g2;
            g4 <= g3;
            
            b1 <= bin;
            b2 <= b1;
            b3 <= b2;
            b4 <= b3;
            
            --Control Signals
            de1 <= de_in;
            de2 <= de1;
            de3 <= de2;
            de4 <= de3;
            
            hs1 <= hs_in;
            hs2 <= hs1;
            hs3 <= hs2;
            hs4 <= hs3;
            
            vs1 <= vs_in;
            vs2 <= vs1;
            vs3 <= vs2;
            vs4 <= vs3;            
            
        end if;
    end process;
    
    
    --Instantiate components
    --TDMS ENCODERS
    r_encoder : tdmi_transmitter port map(
                clk => artificial_base_clk,
                en => artificial_clk_en,
           
                --HDMI Control signals
                CTL => r_ctl,
                DE => de4,
           
                --Data input
                dc => r4,
           
                --Serial Data output output
                TDMI_output => r_tdms_bus    
    );
    
    g_encoder : tdmi_transmitter port map(
                clk => artificial_base_clk,
                en => artificial_clk_en,
           
                --HDMI Control signals
                CTL => g_ctl,
                DE => de4,
           
                --Data input
                dc => g4,
           
                --Serial Data output output
                TDMI_output => g_tdms_bus       
    );
    
    b_encoder : tdmi_transmitter port map(
                clk => artificial_base_clk,
                en => artificial_clk_en,
           
                --HDMI Control signals
                CTL => b_ctl,
                DE => de4,
           
                --Data input
                dc => b4,
           
                --Serial Data output output
                TDMI_output => b_tdms_bus       
    ); 
    
    --SERIALIZERS
    tmds_serialization : tdms_serializer_combined port map(
        data_red => r_tdms_bus,
        data_green => g_tdms_bus,
        data_blue => b_tdms_bus,
        clk => serializer_bit_clk,
        
        --Blue is 0, Green is 1, Red is 2
        TDMS_out => TMDS_stream,
        TDMS_out_not => TMDS_stream_not,
        new_character_clock => TDMS_character_clock,
        en => artificial_clk_en      
    );
    
    --clock generator
    clock_generator : DVI_Clock_Generator port map(
        reset => '0',
        base_clk => clk,
        out_clk_base => artificial_base_clk,
        out_clk_serializer => serializer_bit_clk,
        out_clk_en => artificial_clk_en
    );

end Behavioral;
